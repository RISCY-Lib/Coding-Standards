// The following module does: something
module something (...);

  localparam int SOME_MAGIC_NUMER = 10; // MAGIC_NUMBER is from ...

  ////////////////////
  // Controller FSM //
  ////////////////////
  ...

  ///////////////
  // Data Path //
  ///////////////
  ...

endmodule