if (a == 1'b1) begin
  q <= '0;
end
else begin
  q <= d;
end