always_ff @(posedge clk)
  q <= d;