assign reg_val=((addr==reg_addr)&&enabled)?reg_r:~reg_r;