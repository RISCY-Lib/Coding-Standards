always_ff @(posedge clk) begin
  q <= d;
end