logic [7:0] reg04; // Does not provide any context about what this signal DOES
logic [7:0] status_reg; // Re-made to make the context clearer